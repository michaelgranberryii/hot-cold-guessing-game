library ieee;
use ieee.std_logic_1164.all;

entity debounce_tb is
end debounce_tb;

architecture Behavioral of debounce_tb is

begin

end Behavioral;