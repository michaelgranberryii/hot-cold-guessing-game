library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity number_guess_tb is

end number_guess_tb;

architecture Behavioral of number_guess_tb is

begin

end Behavioral;