library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity single_pulse_detector_tb is

end single_pulse_detector_tb;

architecture Behavioral of single_pulse_detector_tb is

begin

end Behavioral;